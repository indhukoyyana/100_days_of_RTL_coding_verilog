module full_adder(a,b,c,sum,carry);
input a,b,c;
output sum,carry;
assign sum=a^b^c;
assign = (A & B) | (B & Cin) | (A & Cin);
endmodule
